library verilog;
use verilog.vl_types.all;
entity simpleCPU_vlg_vec_tst is
end simpleCPU_vlg_vec_tst;
